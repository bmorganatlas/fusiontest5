["Est exercitationem at ea consequuntur. Rerum nulla soluta et. Consectetur officia distinctio consequatur. Maiores in quas sequi rerum laboriosam.", "Quae maxime nesciunt eius occaecati perspiciatis. Sint aspernatur rerum qui dolorem suscipit. Aliquam ullam odio debitis."]