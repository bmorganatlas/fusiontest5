["Consequatur doloribus odit temporibus hic impedit sint sed. Dolores sed eligendi perspiciatis. Ullam nisi possimus amet quo quasi. Commodi veniam nemo inventore. Repudiandae laborum omnis sunt.", "Quasi dolor minus enim dolores voluptatem in dignissimos. Qui dolorum eos sunt ratione cum. Dolor unde illum laborum quia. Accusamus atque qui eaque.", "Corrupti odit quia illo voluptatem. Aut earum et. Enim nihil architecto inventore placeat et. Deserunt eos autem et ad optio. Dolor numquam laborum.", "Animi quidem vitae. Iure id recusandae sed accusantium at voluptas unde. Soluta cum doloremque in tempore perferendis dolores. Impedit cupiditate voluptas aperiam rem aut. Nam fugiat velit.", "Eos voluptatum animi deserunt rerum atque vel consequatur. Aliquid qui enim. Autem pariatur enim consequatur atque sint. Cupiditate sint nesciunt ratione commodi sed temporibus eos."]