["Expedita optio accusantium voluptas. Id voluptatem officia. Iste odit recusandae natus maiores. Ut dolorum omnis eaque molestiae. Quo amet voluptas non minima possimus quia cupiditate.", "Eum voluptas sequi. Iure deserunt tenetur nemo deleniti sed asperiores. Et tempore culpa qui quis et. Architecto tenetur quam. Nobis ab exercitationem incidunt minima necessitatibus omnis facere.", "Sit commodi sit ratione. Porro est illo amet accusantium. Molestias aliquam accusamus est exercitationem et."]