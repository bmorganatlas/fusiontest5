["Provident quia quos quasi laborum. Cumque occaecati possimus dolor tempore voluptate exercitationem. At nisi vel.", "Et optio qui qui. Debitis voluptatem corporis. Earum totam ratione in velit iste.", "Possimus accusamus inventore odit velit. Aut culpa repudiandae. Aliquid vero quia nisi. Aut autem et.", "Eaque dolores consequatur repudiandae ipsam molestias. Sequi inventore minus voluptas. Expedita dolor est voluptas libero tempore. Velit tempora explicabo aut consequatur.", "Et vel repellendus libero quidem exercitationem quas. Et iste quia numquam molestiae suscipit ut. Dignissimos sit non assumenda ut consequatur. Ea est possimus. Aliquid quaerat ratione omnis quasi est omnis facere.", "Exercitationem molestiae omnis. Officiis corrupti quis quaerat praesentium ut minus consequatur. Maxime vel inventore eligendi est aliquid aut. Omnis asperiores distinctio aut vero rerum nam.", "Aut et ut minima autem vel. Occaecati architecto deleniti dolorem placeat et iure voluptatem. Illo totam id consequuntur ut. Suscipit quia officiis temporibus. Nemo numquam voluptas sint.", "Error quia quas sint consequatur. Distinctio aspernatur exercitationem omnis minus quia vel molestiae. Vel aut maiores. Incidunt tempora aliquid ea alias vero voluptatem labore. Ut inventore expedita dolores.", "Autem ut sint magni. Voluptas eos enim expedita optio vel. Natus in unde veritatis ut cum fuga est. Dolores ut nemo adipisci accusamus voluptas quisquam maiores. Modi consequuntur autem doloremque."]