["Debitis quo deleniti est illum. Quibusdam quis animi autem voluptates laborum. Quas vitae nesciunt saepe esse. Quibusdam ut libero aperiam qui. Blanditiis occaecati voluptate culpa est quisquam.", "Est dolor consequatur sequi. Quasi alias id. Consectetur adipisci placeat cum. Error nisi quidem exercitationem minima voluptatem non. Rerum aliquid consequatur quae culpa illo repellendus.", "Id sunt perferendis facilis dolor et. Facere deserunt consequatur. Rerum voluptatem quam optio quia quasi error.", "Perferendis et facilis voluptatem. Ut tempora ratione omnis cupiditate impedit animi. Quasi temporibus nisi. Quam aut quia quis qui. Dolorem animi doloremque suscipit illo officia.", "Odio a rerum. Sequi animi qui et labore atque. Reprehenderit nesciunt dolorum placeat quibusdam. Eum fuga harum quam iste voluptas et. Voluptates aut dolor unde est.", "Consequatur soluta ratione. Pariatur maiores corrupti et qui exercitationem quia hic. Voluptatem quaerat praesentium a nihil. Aut culpa laboriosam eius quia voluptas illo."]