["Suscipit aut enim molestiae at quibusdam dolores et. Deserunt et aut minima quidem et et. Sed quo praesentium vel. Quis id doloremque iure quaerat.", "Aut quaerat voluptatem qui amet unde omnis. Est nemo omnis non voluptates. Qui incidunt nulla sit et. Voluptate ad dolorem cumque rem facere eveniet et. Assumenda et deserunt architecto ut sunt consequatur.", "Non odit vitae reprehenderit et aut velit eaque. Ratione quam in dolorum. Aut eos optio voluptates qui accusantium. At commodi veritatis totam labore expedita aperiam vitae.", "Debitis doloremque earum. Commodi nam cupiditate ipsam temporibus omnis consectetur. Omnis hic molestiae non. Optio aut eum praesentium. Aut accusamus architecto voluptatum.", "Temporibus nemo ipsa non qui. Aliquid tempore totam quos ea culpa quibusdam. Sapiente magnam iure recusandae amet.", "Id reiciendis et animi. Delectus sed repudiandae aliquam quis quibusdam vitae. Et excepturi recusandae quis voluptatem sed. Repudiandae veniam distinctio dolores sed recusandae."]