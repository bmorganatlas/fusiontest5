["Id earum perspiciatis iure a dicta aut. Saepe cupiditate a earum nemo et similique. Laudantium et qui occaecati. Ut qui labore cumque ducimus culpa consectetur.", "Aut cum molestiae. Et qui sequi odit iste error in. Est eos tenetur illo at unde eveniet. At voluptatem nostrum laudantium sunt.", "Aut numquam perferendis modi quis est. Accusantium aut vero porro accusamus. Minima dolores sint."]