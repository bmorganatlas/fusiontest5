["Est laboriosam natus. Earum laboriosam deleniti et assumenda et non veritatis. Ex nisi ut repellendus id quia. Ab repudiandae consequatur voluptatibus illum voluptas. Cupiditate rem molestiae quam et nostrum.", "Vitae ipsa ex mollitia nesciunt dolor. Harum impedit consectetur. Dolorum qui aut voluptate. Non quia velit et provident optio et aliquid.", "Rerum voluptas repellendus quae est ullam voluptas. Quisquam dolorem eveniet debitis distinctio explicabo. Qui voluptate est.", "Repudiandae quo et. Itaque ipsum quas rem et dicta. Et reiciendis vel molestias voluptate est enim velit. Mollitia quasi aut voluptatem et.", "Et qui quidem quisquam quis accusantium. Dolore repudiandae veniam quia quas aut sed officia. Magnam voluptatem eos placeat. Voluptatem autem quam odio. Ab suscipit odio omnis necessitatibus exercitationem ratione.", "Nisi tenetur vero aut. Et perferendis tempore dolorum dolorem nam et. Praesentium est nemo atque fuga.", "Maiores minima itaque modi sint aut praesentium laborum. Non ut quis consectetur a et. Maxime eligendi est. Dolorem voluptatem asperiores omnis doloremque architecto."]