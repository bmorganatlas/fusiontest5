["Eum et aspernatur animi molestias voluptas recusandae consequatur. Perspiciatis dolorem fugit natus molestias aut vel ipsum. Doloribus nulla corporis reprehenderit dolore maiores dolores.", "Quis aliquid doloribus amet expedita impedit temporibus. Et in sit impedit quis hic. Totam quia culpa optio.", "Sunt vel quasi reiciendis. Molestias exercitationem voluptatibus culpa hic qui vitae quasi. Sed veritatis atque deleniti et ut. Aut quia quod ea qui minus dolorem.", "Qui est veniam nam consequuntur error in totam. Dolorum et pariatur aperiam nostrum libero dolor. A qui voluptatum modi autem voluptatibus facilis. Eveniet doloribus est fugit.", "Aut natus omnis eligendi. Voluptate quia et accusamus. Sint et architecto."]