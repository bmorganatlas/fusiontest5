["Velit rem adipisci harum voluptas dolor. Eos illum saepe sed sit quaerat libero. Ducimus odit excepturi sunt amet ut.", "Asperiores voluptatum voluptas culpa quisquam aut. Quo adipisci non corporis ipsam asperiores velit et. Nobis in soluta. Eaque vitae at laudantium dolores. Dignissimos ipsum ad recusandae et sit est.", "Aut eligendi dolores aliquid. Deleniti doloremque omnis mollitia temporibus ut aut est. Corrupti pariatur similique consequuntur voluptatem qui. Sit tempora consectetur nostrum ad aut quis sapiente. Quia quia quo error."]