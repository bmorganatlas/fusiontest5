["Sint quis voluptates. Rerum iusto expedita voluptas quo. Dolorem vel explicabo velit quisquam cumque.", "Fuga sunt ullam. Doloremque et modi cupiditate nemo minima neque. Quos cupiditate deserunt.", "Aliquid eius nobis magnam. Unde modi qui voluptas labore. Rerum impedit inventore quos sunt. Et nulla est sint nisi.", "Beatae dolorem numquam dicta qui quos deleniti maxime. Est voluptatibus rerum eaque ratione omnis. Magnam nostrum voluptatum illo hic modi.", "Quia aut dolorum iste eveniet vel reprehenderit suscipit. Cupiditate maxime autem ut accusamus vitae quod animi. Incidunt aut quae expedita quis doloribus ea libero.", "Rerum saepe veniam. Ut tempora nam aut tenetur. Consequatur tempore fuga rerum ut numquam et. Quasi qui illo cupiditate. Consequatur deserunt voluptatem et voluptatem nihil.", "Dicta voluptatem rerum eum at magnam ut. Id quasi tempora reiciendis aliquid qui quis consequatur. Dolore quisquam quia veritatis rerum nesciunt. Occaecati magnam animi ipsa sint consequatur iste iure. Dolore vel commodi aliquam."]