["Repudiandae pariatur vel modi. Quidem excepturi voluptates. Velit aut unde sint autem. Consequuntur rerum in minus molestias rerum vel consequatur. Officia consequatur ratione qui sit aspernatur.", "Quasi nesciunt aut omnis modi impedit. Qui et eligendi facilis id dignissimos. Quas ullam itaque exercitationem ipsa ipsum sint et. Pariatur odio dolorum id esse molestiae saepe.", "Est modi veritatis. Rem ducimus debitis qui beatae et dolor. Nostrum est laborum rem et ea. Voluptatem ad labore quasi.", "Voluptatem quae fugiat ipsum quia adipisci magni. Tenetur molestiae et reprehenderit provident magnam explicabo quam. Ut et sapiente tenetur. Quis quia culpa velit. Molestiae autem ex ipsum temporibus."]