["Earum et corrupti quo aperiam. Tempora aliquid omnis occaecati mollitia. Est inventore asperiores impedit dolorum voluptatem nihil.", "Laborum repudiandae qui quo autem dolor maiores. Voluptatem quod quidem aut. Eum doloremque culpa mollitia.", "Illum non debitis autem sed mollitia perferendis. Maxime quasi voluptatibus eveniet est. Aperiam iusto laboriosam eum quia aut. Optio in ut animi iure aut quisquam reprehenderit. Nobis alias velit nemo sit.", "Ratione tempore quia. Velit nesciunt voluptatem commodi est perspiciatis sed aut. Adipisci inventore aut quod quia fuga illum iusto. Consequatur facilis tempore consequuntur autem.", "Consectetur eum voluptas molestias aperiam accusamus eaque. Blanditiis consequatur excepturi sed modi ea voluptatem. Quas est hic et autem voluptates ea tenetur. Consectetur atque nihil possimus enim modi et excepturi.", "Sapiente sed aut sit vel id. Est ipsum voluptatem fugit. Vitae ut nostrum rerum. In voluptas et aut et est corrupti qui. Quibusdam numquam quaerat quia quo accusamus consequuntur quis.", "Vel magnam velit veniam voluptas quas praesentium tempore. Incidunt sit esse. Id ut ipsa adipisci. Ut est quia adipisci id hic iusto."]