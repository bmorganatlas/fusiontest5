["Ad quasi veniam repudiandae cum. Corporis ipsa ut iusto sed dicta et voluptas. Sed dolor nihil placeat cupiditate.", "Est fuga laborum in magni optio sunt rerum. Praesentium odio corporis. Nemo quae eos sapiente.", "Deserunt quia tempore optio aut. Velit sit numquam autem adipisci modi. Officiis atque eaque quis maxime."]