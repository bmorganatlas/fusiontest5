["Sunt at aut. Iusto ut similique facere. Et aspernatur ut velit maxime. Maiores at quia eaque unde tempora.", "Repudiandae sed laboriosam dolorum est aspernatur quas totam. Dignissimos deserunt voluptas ducimus. Soluta est quia consequuntur doloribus. Occaecati laborum recusandae quaerat harum quas. Alias praesentium voluptatem vitae qui sequi."]