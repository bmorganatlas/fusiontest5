["Tempora eius debitis reiciendis dolorum beatae aut. Et voluptate incidunt pariatur alias cupiditate laboriosam. Sed dolorem atque quibusdam dolores. Explicabo sed ea quo dolorum. Fugit enim asperiores temporibus similique aspernatur quia.", "Eius non ex voluptas doloremque. Eos tenetur sequi enim magnam veritatis quo et. Architecto molestiae provident id aliquam quaerat necessitatibus impedit. Eius fugiat est doloremque.", "Voluptas nemo doloribus vel animi. Magnam dignissimos et. A sed quia. Voluptatum eum in.", "Soluta voluptas asperiores. Qui facere facilis ut vel voluptates vitae ad. Aut voluptas debitis illum minus ut ut. Et amet non quis voluptatem quaerat sit ea.", "Corporis aut nesciunt in debitis porro. Et tenetur voluptate voluptates et. Reiciendis aut aut sequi ea veniam deserunt. Veniam cupiditate asperiores error voluptatum.", "Veritatis officia eum sit suscipit cum illum. Rem occaecati distinctio facilis numquam. Explicabo autem ipsum sunt laborum voluptas aliquid. Minus cumque deserunt reprehenderit expedita sed.", "Alias repellendus autem labore. Numquam inventore cum reiciendis libero atque sequi. Blanditiis fugit quas quam rerum nesciunt voluptas. Laudantium veniam nemo itaque excepturi et vero.", "Eligendi ipsam ratione esse quia. Est sint quo sit amet placeat soluta sit. Molestiae laboriosam nisi laudantium consequatur voluptates. Labore exercitationem illum.", "Soluta dolor aspernatur impedit quia. Sit quia autem molestiae dolorem cumque est. Omnis tempore quae. Perferendis quae doloribus quia. Sit in et enim facilis esse."]