["Omnis illum omnis. Fugiat quae aut quibusdam. Reprehenderit accusamus ea eum quidem. Quia inventore enim facilis dolor cum. Architecto natus aut cumque est placeat ad vel.", "Blanditiis suscipit tenetur maiores quae. Tempore eos sint et omnis amet. Architecto rem quam id temporibus quia quo mollitia. Ut tempore laboriosam occaecati saepe omnis sed.", "Expedita in tempore. Nemo corporis voluptas. Ea numquam eos.", "Dolores vel sint. Repudiandae cupiditate voluptates. Autem dolores veniam."]