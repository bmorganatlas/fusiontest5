["Sunt saepe architecto. Dolor eveniet saepe ex et omnis non eum. Ipsum aliquam facilis sequi voluptates inventore at et.", "Reprehenderit est nisi repudiandae. Et voluptas aperiam. Alias ea ratione fugiat laudantium. Tenetur rerum odio quis dolorem repellendus.", "Reprehenderit dolore harum tempore a nesciunt reiciendis. Facilis eius accusantium. Dolor omnis odio.", "Omnis enim rerum quas qui ipsam voluptates dolore. Quia officiis corrupti voluptates tempore. Consequuntur voluptatem blanditiis eos reiciendis temporibus. Consequuntur et deleniti excepturi libero earum facilis.", "Molestiae rem laboriosam temporibus. Est nesciunt ipsam eum odio quia non. Ea omnis sed aut quia perferendis quo rerum. Delectus qui consequatur ut."]