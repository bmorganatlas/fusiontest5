["Totam neque sed et voluptatem nobis temporibus. Veritatis nihil nostrum ullam. Quasi rerum illum saepe.", "Adipisci facilis illo qui perferendis impedit exercitationem voluptas. Blanditiis tempore recusandae et accusantium. Incidunt officia aliquid et. Nesciunt non tenetur illum est ipsum aut.", "Quo quae exercitationem suscipit dolor. Itaque corrupti harum quidem eveniet dolore ullam. Minus labore iste rem omnis. Laudantium in est et quibusdam nam.", "Aliquid ea corporis at fuga. Earum aut eos eligendi. Et error excepturi ut perferendis. Consequuntur eligendi non quis aut ipsa et."]