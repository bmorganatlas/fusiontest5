["Voluptatem quia et consectetur et hic qui et. Itaque iure autem nemo quos. Dolor ea temporibus. Incidunt magnam accusamus aut ad officia.", "Distinctio rem quia eaque natus libero sit qui. Ad quia quam accusantium. Reiciendis asperiores blanditiis aut numquam sed labore.", "Consequatur est vel aliquam. Tempora aut libero. Doloremque qui nihil nihil minus omnis autem.", "Est commodi dolore sint sit. Corporis asperiores minima culpa aut eos velit aliquid. Provident molestias asperiores dolorum aut. Omnis ipsam quis.", "Rerum et in a perspiciatis nemo et. Architecto vitae sit. Non voluptas in et.", "Et nihil minus voluptatem quis alias repellendus est. Saepe ullam dolore dicta tempora. Veniam consequuntur ad nam aut porro. Distinctio odio ea ipsam. Eligendi qui et praesentium.", "Laudantium quia omnis molestias. Iusto nihil reiciendis rem explicabo. Ad minus deserunt."]