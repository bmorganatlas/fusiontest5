["Officiis veritatis sit. Est aut voluptatem sequi. Tempora earum magni eius impedit rerum. Eius neque odio voluptatibus eum.", "Vel et velit voluptate. Ipsam enim incidunt placeat perferendis quos. Deserunt tempora est.", "Sed dolorum laborum dicta optio ut alias reiciendis. Aliquid sit inventore laboriosam rerum. Ipsum deleniti odio et rerum.", "Vitae sit aut aut rerum. Sit magni voluptatem. Ipsa assumenda architecto rem omnis voluptas labore ducimus.", "Voluptatum nesciunt tenetur aut error magnam unde. Dolor labore debitis earum. Fugit aliquam optio. Voluptatem quia doloribus voluptas.", "Aliquid doloremque beatae laborum. Aut recusandae et et. Soluta rem autem ipsa sint.", "Inventore quia similique reprehenderit officiis aut. Est repudiandae harum. Perspiciatis enim explicabo culpa alias neque consectetur provident.", "Rerum dolore qui. Voluptatem excepturi debitis aperiam magnam soluta. Provident non a exercitationem. Est explicabo tempore optio omnis iste recusandae.", "Sed saepe et. Modi eveniet dolor ex tenetur sit animi. Alias ut vel. Culpa repellat eaque architecto aut nostrum.", "Suscipit voluptas est est et. Ratione nesciunt quia omnis harum recusandae. Adipisci suscipit et quas recusandae."]