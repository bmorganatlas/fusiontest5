["Atque nam omnis aut. Est eos qui odio voluptatem. Culpa nam porro quos. Praesentium magnam fuga autem soluta. A doloribus modi eveniet sit pariatur praesentium fugit.", "Non commodi et quis qui saepe facere. Eum ut commodi ea. Nam animi et id commodi cum.", "Quas error id culpa harum corrupti cumque exercitationem. Sunt quam doloremque. Voluptatem et autem corporis ut deleniti sapiente inventore.", "Est reprehenderit id amet. Rem aspernatur eligendi et. Quis non cumque. Corrupti et sed.", "Ut amet adipisci voluptatem voluptatem reiciendis quam. Voluptas deleniti saepe doloribus qui velit veritatis. Delectus dolor minus quia accusantium voluptas. Doloribus rerum iusto harum. Nihil rerum ratione laudantium similique.", "Voluptatem consequatur cumque distinctio aspernatur iusto. Voluptas nihil et laudantium rerum quo nulla. Molestias consectetur dolores.", "Autem eaque est voluptas reiciendis quia dicta. Rem adipisci eaque qui possimus deleniti praesentium sint. Aut id veritatis sit suscipit.", "Atque illo enim. Dicta ad et ex placeat qui culpa. A praesentium quia. Commodi at facilis laborum architecto molestiae.", "Incidunt soluta est ipsam. Qui eum tempore. Itaque nemo labore sapiente saepe voluptas eaque. Quos unde laudantium aut."]