["Repudiandae beatae dolore qui eveniet. Voluptas quae ab dolorem dolores ut vel atque. Incidunt est nemo totam similique dolorem repellendus corporis. Deleniti veritatis eligendi ipsa voluptatem. Nemo et modi.", "Dolor sed ullam. Voluptates itaque enim non. Aperiam tempore vel. Quis asperiores perspiciatis nihil itaque dolore.", "Sed eaque vel suscipit rerum dignissimos ad et. Qui officiis quibusdam. Impedit fuga illo odit et. Totam eaque et asperiores eum exercitationem sed illo."]