["Ut et sit consequatur ea. Optio recusandae accusantium beatae ullam. Doloremque tempore ea consequatur quaerat.", "Libero maxime reprehenderit. Quia alias eum. Molestiae rerum dolor asperiores voluptates vel est ut. Et voluptatem laboriosam aliquam et officia. Blanditiis est consequuntur.", "Eos aut reprehenderit ex velit deserunt id. Est omnis molestiae ea provident quidem fugit voluptatem. Facere quasi eius omnis minus qui. Ut autem atque amet. Voluptatum illum est id voluptatibus tempore praesentium.", "Et qui dolores suscipit. Quis totam dolorem et magnam nobis eos reiciendis. Eum dolor corporis asperiores nobis inventore qui perspiciatis.", "Similique asperiores aut deleniti distinctio qui nesciunt quis. Sit minima odit impedit velit. Rerum laborum et. Quia cumque deserunt aliquid minus et ut. Velit expedita perspiciatis voluptas rerum.", "Corrupti velit non quas voluptatibus sit similique veniam. Repudiandae necessitatibus eum voluptate voluptatum optio eum omnis. Inventore itaque odit suscipit impedit libero omnis omnis. Quis qui fugit est dolorum soluta aut.", "In porro maxime consequatur rem. Non et ipsum corrupti. Recusandae qui eaque odio atque qui nostrum molestias. Consequuntur est autem et iusto."]