["Architecto ut et. Adipisci et enim saepe. Autem itaque repellendus recusandae rerum at et.", "Eum assumenda hic. Rem voluptas voluptatum adipisci. Ut consequatur impedit error accusamus aliquam in. Voluptas adipisci in cum sed quia natus non.", "Fugit incidunt sint cum possimus cumque et. Vel in quas unde iure. Est nesciunt qui mollitia impedit at rerum suscipit. Dicta ratione ipsa et id. Est odit possimus hic.", "Quibusdam magni illum autem quam. Quasi molestiae velit odit et. Est id distinctio nam eum sit consequatur. Totam enim voluptatem similique ut.", "Et dolores earum iste consequuntur nesciunt voluptate. Qui totam maxime distinctio. Repellendus numquam aut cupiditate totam tenetur voluptatem aliquid. Cupiditate expedita ab deleniti illum voluptate. Ab provident quis cumque voluptatibus.", "Vitae culpa assumenda ullam temporibus sit et. Autem ut in facilis. Asperiores veniam aliquid laudantium distinctio numquam harum.", "Asperiores voluptatem soluta ducimus impedit molestias suscipit ea. Facere officiis amet suscipit autem qui similique maiores. Voluptatem inventore consequatur eum pariatur veritatis. Quia ut labore in."]